// Naive Implementation of Linear Layer using Rotation Algorithm
module linear_layer (
    input [63:0] x0, x1, x2, x3, x4,
    output [63:0] o0, o1, o2, o3, o4
);

    assign o0 = x0 ^ ((x0 >> 19) | ((x0 & (1<<19)-1) << (64-19))) ^ ((x0 >> 28) | ((x0 & (1<<28)-1) << (64-28)));
    assign o1 = x1 ^ ((x1 >> 61) | ((x1 & (1<<61)-1) << (64-61))) ^ ((x1 >> 39) | ((x1 & (1<<39)-1) << (64-39)));
    assign o2 = x2 ^ ((x2 >> 1)  | ((x2 & (1<<1)-1) << (64-1)))   ^ ((x2 >> 6)  | ((x2 & (1<<6)-1)  << (64-6)));
    assign o3 = x3 ^ ((x3 >> 10) | ((x3 & (1<<10)-1) << (64-10))) ^ ((x3 >> 17) | ((x3 & (1<<17)-1) << (64-17)));
    assign o4 = x4 ^ ((x4 >> 7)  | ((x4 & (1<<7)-1) << (64-7)))   ^ ((x4 >> 41) | ((x4 & (1<<41)-1) << (64-41)));
endmodule