// Optimized Linear Layer using Matrix Multiplication Algorithm
module linear_layer (
    input [63:0] X0, X1, X2, X3, X4,
    output [63:0] Y0, Y1, Y2, Y3, Y4
);
    wire [319:0] s;
    assign s = {X0, X1, X2, X3, X4};

    assign Y0 = {(s[319] ^ s[283] ^ s[274]), (s[318] ^ s[282] ^ s[273]), (s[317] ^ s[281] ^ s[272]), (s[316] ^ s[280] ^ s[271]), (s[315] ^ s[279] ^ s[270]), (s[314] ^ s[278] ^ s[269]), (s[313] ^ s[277] ^ s[268]), (s[312] ^ s[276] ^ s[267]),
                (s[311] ^ s[275] ^ s[266]), (s[310] ^ s[274] ^ s[265]), (s[309] ^ s[273] ^ s[264]), (s[308] ^ s[272] ^ s[263]), (s[307] ^ s[271] ^ s[262]), (s[306] ^ s[270] ^ s[261]), (s[305] ^ s[269] ^ s[260]), (s[304] ^ s[268] ^ s[259]),
                (s[303] ^ s[267] ^ s[258]), (s[302] ^ s[266] ^ s[257]), (s[301] ^ s[265] ^ s[256]), (s[319] ^ s[300] ^ s[264]), (s[318] ^ s[299] ^ s[263]), (s[317] ^ s[298] ^ s[262]), (s[316] ^ s[297] ^ s[261]), (s[315] ^ s[296] ^ s[260]),
                (s[314] ^ s[295] ^ s[259]), (s[313] ^ s[294] ^ s[258]), (s[312] ^ s[293] ^ s[257]), (s[311] ^ s[292] ^ s[256]), (s[319] ^ s[310] ^ s[291]), (s[318] ^ s[309] ^ s[290]), (s[317] ^ s[308] ^ s[289]), (s[316] ^ s[307] ^ s[288]),
                (s[315] ^ s[306] ^ s[287]), (s[314] ^ s[305] ^ s[286]), (s[313] ^ s[304] ^ s[285]), (s[312] ^ s[303] ^ s[284]), (s[311] ^ s[302] ^ s[283]), (s[310] ^ s[301] ^ s[282]), (s[309] ^ s[300] ^ s[281]), (s[308] ^ s[299] ^ s[280]),
                (s[307] ^ s[298] ^ s[279]), (s[306] ^ s[297] ^ s[278]), (s[305] ^ s[296] ^ s[277]), (s[304] ^ s[295] ^ s[276]), (s[303] ^ s[294] ^ s[275]), (s[302] ^ s[293] ^ s[274]), (s[301] ^ s[292] ^ s[273]), (s[300] ^ s[291] ^ s[272]),
                (s[299] ^ s[290] ^ s[271]), (s[298] ^ s[289] ^ s[270]), (s[297] ^ s[288] ^ s[269]), (s[296] ^ s[287] ^ s[268]), (s[295] ^ s[286] ^ s[267]), (s[294] ^ s[285] ^ s[266]), (s[293] ^ s[284] ^ s[265]), (s[292] ^ s[283] ^ s[264]),
                (s[291] ^ s[282] ^ s[263]), (s[290] ^ s[281] ^ s[262]), (s[289] ^ s[280] ^ s[261]), (s[288] ^ s[279] ^ s[260]), (s[287] ^ s[278] ^ s[259]), (s[286] ^ s[277] ^ s[258]), (s[285] ^ s[276] ^ s[257]), (s[284] ^ s[275] ^ s[256])};

    assign Y1 = {(s[255] ^ s[252] ^ s[230]), (s[254] ^ s[251] ^ s[229]), (s[253] ^ s[250] ^ s[228]), (s[252] ^ s[249] ^ s[227]), (s[251] ^ s[248] ^ s[226]), (s[250] ^ s[247] ^ s[225]), (s[249] ^ s[246] ^ s[224]), (s[248] ^ s[245] ^ s[223]),
                (s[247] ^ s[244] ^ s[222]), (s[246] ^ s[243] ^ s[221]), (s[245] ^ s[242] ^ s[220]), (s[244] ^ s[241] ^ s[219]), (s[243] ^ s[240] ^ s[218]), (s[242] ^ s[239] ^ s[217]), (s[241] ^ s[238] ^ s[216]), (s[240] ^ s[237] ^ s[215]),
                (s[239] ^ s[236] ^ s[214]), (s[238] ^ s[235] ^ s[213]), (s[237] ^ s[234] ^ s[212]), (s[236] ^ s[233] ^ s[211]), (s[235] ^ s[232] ^ s[210]), (s[234] ^ s[231] ^ s[209]), (s[233] ^ s[230] ^ s[208]), (s[232] ^ s[229] ^ s[207]),
                (s[231] ^ s[228] ^ s[206]), (s[230] ^ s[227] ^ s[205]), (s[229] ^ s[226] ^ s[204]), (s[228] ^ s[225] ^ s[203]), (s[227] ^ s[224] ^ s[202]), (s[226] ^ s[223] ^ s[201]), (s[225] ^ s[222] ^ s[200]), (s[224] ^ s[221] ^ s[199]),
                (s[223] ^ s[220] ^ s[198]), (s[222] ^ s[219] ^ s[197]), (s[221] ^ s[218] ^ s[196]), (s[220] ^ s[217] ^ s[195]), (s[219] ^ s[216] ^ s[194]), (s[218] ^ s[215] ^ s[193]), (s[217] ^ s[214] ^ s[192]), (s[255] ^ s[216] ^ s[213]),
                (s[254] ^ s[215] ^ s[212]), (s[253] ^ s[214] ^ s[211]), (s[252] ^ s[213] ^ s[210]), (s[251] ^ s[212] ^ s[209]), (s[250] ^ s[211] ^ s[208]), (s[249] ^ s[210] ^ s[207]), (s[248] ^ s[209] ^ s[206]), (s[247] ^ s[208] ^ s[205]),
                (s[246] ^ s[207] ^ s[204]), (s[245] ^ s[206] ^ s[203]), (s[244] ^ s[205] ^ s[202]), (s[243] ^ s[204] ^ s[201]), (s[242] ^ s[203] ^ s[200]), (s[241] ^ s[202] ^ s[199]), (s[240] ^ s[201] ^ s[198]), (s[239] ^ s[200] ^ s[197]),
                (s[238] ^ s[199] ^ s[196]), (s[237] ^ s[198] ^ s[195]), (s[236] ^ s[197] ^ s[194]), (s[235] ^ s[196] ^ s[193]), (s[234] ^ s[195] ^ s[192]), (s[255] ^ s[233] ^ s[194]), (s[254] ^ s[232] ^ s[193]), (s[253] ^ s[231] ^ s[192])};

    assign Y2 = {(s[191] ^ s[133] ^ s[128]), (s[191] ^ s[190] ^ s[132]), (s[190] ^ s[189] ^ s[131]), (s[189] ^ s[188] ^ s[130]), (s[188] ^ s[187] ^ s[129]), (s[187] ^ s[186] ^ s[128]), (s[191] ^ s[186] ^ s[185]), (s[190] ^ s[185] ^ s[184]),
                (s[189] ^ s[184] ^ s[183]), (s[188] ^ s[183] ^ s[182]), (s[187] ^ s[182] ^ s[181]), (s[186] ^ s[181] ^ s[180]), (s[185] ^ s[180] ^ s[179]), (s[184] ^ s[179] ^ s[178]), (s[183] ^ s[178] ^ s[177]), (s[182] ^ s[177] ^ s[176]),
                (s[181] ^ s[176] ^ s[175]), (s[180] ^ s[175] ^ s[174]), (s[179] ^ s[174] ^ s[173]), (s[178] ^ s[173] ^ s[172]), (s[177] ^ s[172] ^ s[171]), (s[176] ^ s[171] ^ s[170]), (s[175] ^ s[170] ^ s[169]), (s[174] ^ s[169] ^ s[168]),
                (s[173] ^ s[168] ^ s[167]), (s[172] ^ s[167] ^ s[166]), (s[171] ^ s[166] ^ s[165]), (s[170] ^ s[165] ^ s[164]), (s[169] ^ s[164] ^ s[163]), (s[168] ^ s[163] ^ s[162]), (s[167] ^ s[162] ^ s[161]), (s[166] ^ s[161] ^ s[160]),
                (s[165] ^ s[160] ^ s[159]), (s[164] ^ s[159] ^ s[158]), (s[163] ^ s[158] ^ s[157]), (s[162] ^ s[157] ^ s[156]), (s[161] ^ s[156] ^ s[155]), (s[160] ^ s[155] ^ s[154]), (s[159] ^ s[154] ^ s[153]), (s[158] ^ s[153] ^ s[152]),
                (s[157] ^ s[152] ^ s[151]), (s[156] ^ s[151] ^ s[150]), (s[155] ^ s[150] ^ s[149]), (s[154] ^ s[149] ^ s[148]), (s[153] ^ s[148] ^ s[147]), (s[152] ^ s[147] ^ s[146]), (s[151] ^ s[146] ^ s[145]), (s[150] ^ s[145] ^ s[144]),
                (s[149] ^ s[144] ^ s[143]), (s[148] ^ s[143] ^ s[142]), (s[147] ^ s[142] ^ s[141]), (s[146] ^ s[141] ^ s[140]), (s[145] ^ s[140] ^ s[139]), (s[144] ^ s[139] ^ s[138]), (s[143] ^ s[138] ^ s[137]), (s[142] ^ s[137] ^ s[136]),
                (s[141] ^ s[136] ^ s[135]), (s[140] ^ s[135] ^ s[134]), (s[139] ^ s[134] ^ s[133]), (s[138] ^ s[133] ^ s[132]), (s[137] ^ s[132] ^ s[131]), (s[136] ^ s[131] ^ s[130]), (s[135] ^ s[130] ^ s[129]), (s[134] ^ s[129] ^ s[128])};

    assign Y3 = {(s[127] ^ s[80] ^ s[73]), (s[126] ^ s[79] ^ s[72]), (s[125] ^ s[78] ^ s[71]), (s[124] ^ s[77] ^ s[70]), (s[123] ^ s[76] ^ s[69]), (s[122] ^ s[75] ^ s[68]), (s[121] ^ s[74] ^ s[67]), (s[120] ^ s[73] ^ s[66]),
                (s[119] ^ s[72] ^ s[65]), (s[118] ^ s[71] ^ s[64]), (s[127] ^ s[117] ^ s[70]), (s[126] ^ s[116] ^ s[69]), (s[125] ^ s[115] ^ s[68]), (s[124] ^ s[114] ^ s[67]), (s[123] ^ s[113] ^ s[66]), (s[122] ^ s[112] ^ s[65]),
                (s[121] ^ s[111] ^ s[64]), (s[127] ^ s[120] ^ s[110]), (s[126] ^ s[119] ^ s[109]), (s[125] ^ s[118] ^ s[108]), (s[124] ^ s[117] ^ s[107]), (s[123] ^ s[116] ^ s[106]), (s[122] ^ s[115] ^ s[105]), (s[121] ^ s[114] ^ s[104]),
                (s[120] ^ s[113] ^ s[103]), (s[119] ^ s[112] ^ s[102]), (s[118] ^ s[111] ^ s[101]), (s[117] ^ s[110] ^ s[100]), (s[116] ^ s[109] ^ s[99]), (s[115] ^ s[108] ^ s[98]), (s[114] ^ s[107] ^ s[97]), (s[113] ^ s[106] ^ s[96]),
                (s[112] ^ s[105] ^ s[95]), (s[111] ^ s[104] ^ s[94]), (s[110] ^ s[103] ^ s[93]), (s[109] ^ s[102] ^ s[92]), (s[108] ^ s[101] ^ s[91]), (s[107] ^ s[100] ^ s[90]), (s[106] ^ s[99] ^ s[89]), (s[105] ^ s[98] ^ s[88]),
                (s[104] ^ s[97] ^ s[87]), (s[103] ^ s[96] ^ s[86]), (s[102] ^ s[95] ^ s[85]), (s[101] ^ s[94] ^ s[84]), (s[100] ^ s[93] ^ s[83]), (s[99] ^ s[92] ^ s[82]), (s[98] ^ s[91] ^ s[81]), (s[97] ^ s[90] ^ s[80]),
                (s[96] ^ s[89] ^ s[79]), (s[95] ^ s[88] ^ s[78]), (s[94] ^ s[87] ^ s[77]), (s[93] ^ s[86] ^ s[76]), (s[92] ^ s[85] ^ s[75]), (s[91] ^ s[84] ^ s[74]), (s[90] ^ s[83] ^ s[73]), (s[89] ^ s[82] ^ s[72]),
                (s[88] ^ s[81] ^ s[71]), (s[87] ^ s[80] ^ s[70]), (s[86] ^ s[79] ^ s[69]), (s[85] ^ s[78] ^ s[68]), (s[84] ^ s[77] ^ s[67]), (s[83] ^ s[76] ^ s[66]), (s[82] ^ s[75] ^ s[65]), (s[81] ^ s[74] ^ s[64])};

    assign Y4 = {(s[63] ^ s[40] ^ s[6]), (s[62] ^ s[39] ^ s[5]), (s[61] ^ s[38] ^ s[4]), (s[60] ^ s[37] ^ s[3]), (s[59] ^ s[36] ^ s[2]), (s[58] ^ s[35] ^ s[1]), (s[57] ^ s[34] ^ s[0]), (s[63] ^ s[56] ^ s[33]),
                (s[62] ^ s[55] ^ s[32]), (s[61] ^ s[54] ^ s[31]), (s[60] ^ s[53] ^ s[30]), (s[59] ^ s[52] ^ s[29]), (s[58] ^ s[51] ^ s[28]), (s[57] ^ s[50] ^ s[27]), (s[56] ^ s[49] ^ s[26]), (s[55] ^ s[48] ^ s[25]),
                (s[54] ^ s[47] ^ s[24]), (s[53] ^ s[46] ^ s[23]), (s[52] ^ s[45] ^ s[22]), (s[51] ^ s[44] ^ s[21]), (s[50] ^ s[43] ^ s[20]), (s[49] ^ s[42] ^ s[19]), (s[48] ^ s[41] ^ s[18]), (s[47] ^ s[40] ^ s[17]),
                (s[46] ^ s[39] ^ s[16]), (s[45] ^ s[38] ^ s[15]), (s[44] ^ s[37] ^ s[14]), (s[43] ^ s[36] ^ s[13]), (s[42] ^ s[35] ^ s[12]), (s[41] ^ s[34] ^ s[11]), (s[40] ^ s[33] ^ s[10]), (s[39] ^ s[32] ^ s[9]),
                (s[38] ^ s[31] ^ s[8]), (s[37] ^ s[30] ^ s[7]), (s[36] ^ s[29] ^ s[6]), (s[35] ^ s[28] ^ s[5]), (s[34] ^ s[27] ^ s[4]), (s[33] ^ s[26] ^ s[3]), (s[32] ^ s[25] ^ s[2]), (s[31] ^ s[24] ^ s[1]),
                (s[30] ^ s[23] ^ s[0]), (s[63] ^ s[29] ^ s[22]), (s[62] ^ s[28] ^ s[21]), (s[61] ^ s[27] ^ s[20]), (s[60] ^ s[26] ^ s[19]), (s[59] ^ s[25] ^ s[18]), (s[58] ^ s[24] ^ s[17]), (s[57] ^ s[23] ^ s[16]),
                (s[56] ^ s[22] ^ s[15]), (s[55] ^ s[21] ^ s[14]), (s[54] ^ s[20] ^ s[13]), (s[53] ^ s[19] ^ s[12]), (s[52] ^ s[18] ^ s[11]), (s[51] ^ s[17] ^ s[10]), (s[50] ^ s[16] ^ s[9]), (s[49] ^ s[15] ^ s[8]),
                (s[48] ^ s[14] ^ s[7]), (s[47] ^ s[13] ^ s[6]), (s[46] ^ s[12] ^ s[5]), (s[45] ^ s[11] ^ s[4]), (s[44] ^ s[10] ^ s[3]), (s[43] ^ s[9] ^ s[2]), (s[42] ^ s[8] ^ s[1]), (s[41] ^ s[7] ^ s[0])};

endmodule

/*
S[0] = [s0 + s36 + s45, s1 + s37 + s46, s2 + s38 + s47, s3 + s39 + s48, s4 + s40 + s49, s5 + s41 + s50, s6 + s42 + s51, s7 + s43 + s52, s8 + s44 + s53, s9 + s45 + s54, s10 + s46 + s55, s11 + s47 + s56, s12 + s48 + s57, s13 + s49 + s58, s14 + s50 + s59, s15 + s51 + s60, s16 + s52 + s61, s17 + s53 + s62, s18 + s54 + s63, s0 + s19 + s55, s1 + s20 + s56, s2 + s21 + s57, s3 + s22 + s58, s4 + s23 + s59, s5 + s24 + s60, s6 + s25 + s61, s7 + s26 + s62, s8 + s27 + s63, s0 + s9 + s28, s1 + s10 + s29, s2 + s11 + s30, s3 + s12 + s31, s4 + s13 + s32, s5 + s14 + s33, s6 + s15 + s34, s7 + s16 + s35, s8 + s17 + s36, s9 + s18 + s37, s10 + s19 + s38, s11 + s20 + s39, s12 + s21 + s40, s13 + s22 + s41, s14 + s23 + s42, s15 + s24 + s43, s16 + s25 + s44, s17 + s26 + s45, s18 + s27 + s46, s19 + s28 + s47, s20 + s29 + s48, s21 + s30 + s49, s22 + s31 + s50, s23 + s32 + s51, s24 + s33 + s52, s25 + s34 + s53, s26 + s35 + s54, s27 + s36 + s55, s28 + s37 + s56, s29 + s38 + s57, s30 + s39 + s58, s31 + s40 + s59, s32 + s41 + s60, s33 + s42 + s61, s34 + s43 + s62, s35 + s44 + s63]
S[1] = [s64 + s67 + s89, s65 + s68 + s90, s66 + s69 + s91, s67 + s70 + s92, s68 + s71 + s93, s69 + s72 + s94, s70 + s73 + s95, s71 + s74 + s96, s72 + s75 + s97, s73 + s76 + s98, s74 + s77 + s99, s75 + s78 + s100, s76 + s79 + s101, s77 + s80 + s102, s78 + s81 + s103, s79 + s82 + s104, s80 + s83 + s105, s81 + s84 + s106, s82 + s85 + s107, s83 + s86 + s108, s84 + s87 + s109, s85 + s88 + s110, s86 + s89 + s111, s87 + s90 + s112, s88 + s91 + s113, s89 + s92 + s114, s90 + s93 + s115, s91 + s94 + s116, s92 + s95 + s117, s93 + s96 + s118, s94 + s97 + s119, s95 + s98 + s120, s96 + s99 + s121, s97 + s100 + s122, s98 + s101 + s123, s99 + s102 + s124, s100 + s103 + s125, s101 + s104 + s126, s102 + s105 + s127, s64 + s103 + s106, s65 + s104 + s107, s66 + s105 + s108, s67 + s106 + s109, s68 + s107 + s110, s69 + s108 + s111, s70 + s109 + s112, s71 + s110 + s113, s72 + s111 + s114, s73 + s112 + s115, s74 + s113 + s116, s75 + s114 + s117, s76 + s115 + s118, s77 + s116 + s119, s78 + s117 + s120, s79 + s118 + s121, s80 + s119 + s122, s81 + s120 + s123, s82 + s121 + s124, s83 + s122 + s125, s84 + s123 + s126, s85 + s124 + s127, s64 + s86 + s125, s65 + s87 + s126, s66 + s88 + s127]
S[2] = [s128 + s186 + s191, s128 + s129 + s187, s129 + s130 + s188, s130 + s131 + s189, s131 + s132 + s190, s132 + s133 + s191, s128 + s133 + s134, s129 + s134 + s135, s130 + s135 + s136, s131 + s136 + s137, s132 + s137 + s138, s133 + s138 + s139, s134 + s139 + s140, s135 + s140 + s141, s136 + s141 + s142, s137 + s142 + s143, s138 + s143 + s144, s139 + s144 + s145, s140 + s145 + s146, s141 + s146 + s147, s142 + s147 + s148, s143 + s148 + s149, s144 + s149 + s150, s145 + s150 + s151, s146 + s151 + s152, s147 + s152 + s153, s148 + s153 + s154, s149 + s154 + s155, s150 + s155 + s156, s151 + s156 + s157, s152 + s157 + s158, s153 + s158 + s159, s154 + s159 + s160, s155 + s160 + s161, s156 + s161 + s162, s157 + s162 + s163, s158 + s163 + s164, s159 + s164 + s165, s160 + s165 + s166, s161 + s166 + s167, s162 + s167 + s168, s163 + s168 + s169, s164 + s169 + s170, s165 + s170 + s171, s166 + s171 + s172, s167 + s172 + s173, s168 + s173 + s174, s169 + s174 + s175, s170 + s175 + s176, s171 + s176 + s177, s172 + s177 + s178, s173 + s178 + s179, s174 + s179 + s180, s175 + s180 + s181, s176 + s181 + s182, s177 + s182 + s183, s178 + s183 + s184, s179 + s184 + s185, s180 + s185 + s186, s181 + s186 + s187, s182 + s187 + s188, s183 + s188 + s189, s184 + s189 + s190, s185 + s190 + s191]
S[3] = [s192 + s239 + s246, s193 + s240 + s247, s194 + s241 + s248, s195 + s242 + s249, s196 + s243 + s250, s197 + s244 + s251, s198 + s245 + s252, s199 + s246 + s253, s200 + s247 + s254, s201 + s248 + s255, s192 + s202 + s249, s193 + s203 + s250, s194 + s204 + s251, s195 + s205 + s252, s196 + s206 + s253, s197 + s207 + s254, s198 + s208 + s255, s192 + s199 + s209, s193 + s200 + s210, s194 + s201 + s211, s195 + s202 + s212, s196 + s203 + s213, s197 + s204 + s214, s198 + s205 + s215, s199 + s206 + s216, s200 + s207 + s217, s201 + s208 + s218, s202 + s209 + s219, s203 + s210 + s220, s204 + s211 + s221, s205 + s212 + s222, s206 + s213 + s223, s207 + s214 + s224, s208 + s215 + s225, s209 + s216 + s226, s210 + s217 + s227, s211 + s218 + s228, s212 + s219 + s229, s213 + s220 + s230, s214 + s221 + s231, s215 + s222 + s232, s216 + s223 + s233, s217 + s224 + s234, s218 + s225 + s235, s219 + s226 + s236, s220 + s227 + s237, s221 + s228 + s238, s222 + s229 + s239, s223 + s230 + s240, s224 + s231 + s241, s225 + s232 + s242, s226 + s233 + s243, s227 + s234 + s244, s228 + s235 + s245, s229 + s236 + s246, s230 + s237 + s247, s231 + s238 + s248, s232 + s239 + s249, s233 + s240 + s250, s234 + s241 + s251, s235 + s242 + s252, s236 + s243 + s253, s237 + s244 + s254, s238 + s245 + s255]
S[4] = [s256 + s279 + s313, s257 + s280 + s314, s258 + s281 + s315, s259 + s282 + s316, s260 + s283 + s317, s261 + s284 + s318, s262 + s285 + s319, s256 + s263 + s286, s257 + s264 + s287, s258 + s265 + s288, s259 + s266 + s289, s260 + s267 + s290, s261 + s268 + s291, s262 + s269 + s292, s263 + s270 + s293, s264 + s271 + s294, s265 + s272 + s295, s266 + s273 + s296, s267 + s274 + s297, s268 + s275 + s298, s269 + s276 + s299, s270 + s277 + s300, s271 + s278 + s301, s272 + s279 + s302, s273 + s280 + s303, s274 + s281 + s304, s275 + s282 + s305, s276 + s283 + s306, s277 + s284 + s307, s278 + s285 + s308, s279 + s286 + s309, s280 + s287 + s310, s281 + s288 + s311, s282 + s289 + s312, s283 + s290 + s313, s284 + s291 + s314, s285 + s292 + s315, s286 + s293 + s316, s287 + s294 + s317, s288 + s295 + s318, s289 + s296 + s319, s256 + s290 + s297, s257 + s291 + s298, s258 + s292 + s299, s259 + s293 + s300, s260 + s294 + s301, s261 + s295 + s302, s262 + s296 + s303, s263 + s297 + s304, s264 + s298 + s305, s265 + s299 + s306, s266 + s300 + s307, s267 + s301 + s308, s268 + s302 + s309, s269 + s303 + s310, s270 + s304 + s311, s271 + s305 + s312, s272 + s306 + s313, s273 + s307 + s314, s274 + s308 + s315, s275 + s309 + s316, s276 + s310 + s317, s277 + s311 + s318, s278 + s312 + s319]
*/