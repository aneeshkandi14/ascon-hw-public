module sub_layer_ti (
    input x0_0,x1_0,x2_0,x3_0,x4_0,
    input x0_1,x1_1,x2_1,x3_1,x4_1,
    input x0_2,x1_2,x2_2,x3_2,x4_2,

    output y0_0,y1_0,y2_0,y3_0,y4_0
);

    assign y0_0 = (x4_0 & x1_0) ^ (x4_0 & x1_2) ^ (x4_2 & x1_0) ^ x3_2 ^ (x2_0 & x1_2) ^ (x2_2 & x1_0) ^ x2_2 ^ (x1_0 & x0_2) ^ x1_0 ^ (x1_2 & x0_0) ^ (x1_2 & x0_2) ;
    assign y1_0 = x4_1 ^ (x3_1 & x2_1) ^ (x3_1 & x2_2) ^ (x3_1 & x1_2) ^ x3_1 ^ (x3_2 & x2_1) ^ (x3_2 & x1_1) ^ (x3_2 & x1_2) ^ x3_2 ^ (x2_1 & x1_2) ^ x2_1 ^ (x2_2 & x1_1) ^ (x2_2 & x1_2) ^ x0_1 ^ x0_2 ;
    assign y2_0 = (x4_0 & x3_0) ^ (x4_0 & x3_2) ^ x4_0 ^ (x4_2 & x3_0) ^ (x4_2 & x3_2) ^ x2_2 ^ x1_0 ;
    assign y3_0 = (x4_1 & x0_2) ^ x4_1 ^ (x4_2 & x0_1) ^ x4_2 ^ (x3_1 & x0_1) ^ (x3_1 & x0_2) ^ (x3_2 & x0_1) ^ (x3_2 & x0_2) ^ x2_1 ^ x1_2 ;
    assign y4_0 = (x4_1 & x1_2) ^ (x4_2 & x1_1) ^ x3_1 ^ (x1_1 & x0_1) ^ (x1_1 & x0_2) ^ (x1_2 & x0_1) ^ x1_2 ;

    assign y0_1 = (x4_0 & x1_1) ^ (x4_1 & x1_0) ^ (x4_1 & x1_1) ^ x3_0 ^ (x2_0 & x1_0) ^ (x2_0 & x1_1) ^ x2_0 ^ (x2_1 & x1_0) ^ x2_1 ^ (x1_0 & x0_0) ^ (x1_0 & x0_1) ^ (x1_1 & x0_0) ^ x1_1 ^ x0_0 ^ x0_1 ;
    assign y1_1 = x4_0 ^ (x3_0 & x2_0) ^ (x3_0 & x2_1) ^ (x3_0 & x1_0) ^ (x3_0 & x1_1) ^ x3_0 ^ (x3_1 & x2_0) ^ (x3_1 & x1_0) ^ (x3_1 & x1_1) ^ (x2_0 & x1_1) ^ (x2_1 & x1_0) ^ (x2_1 & x1_1) ^ x1_1 ^ x0_0 ;
    assign y2_1 = (x4_1 & x3_1) ^ (x4_1 & x3_2) ^ x4_1 ^ (x4_2 & x3_1) ^ x4_2 ^ x2_1 ^ x1_2 ;
    assign y3_1 = (x4_0 & x0_0) ^ (x4_0 & x0_1) ^ x4_0 ^ (x4_1 & x0_0) ^ (x4_1 & x0_1) ^ (x3_0 & x0_0) ^ (x3_0 & x0_1) ^ x3_0 ^ (x3_1 & x0_0) ^ x3_1 ^ x2_0 ^ x1_1 ^ x0_1 ;
    assign y4_1 = (x4_0 & x1_1) ^ x4_0 ^ (x4_1 & x1_0) ^ (x4_1 & x1_1) ^ x4_1 ^ (x1_0 & x0_0) ^ (x1_0 & x0_1) ^ x1_0 ^ (x1_1 & x0_0) ^ x1_1 ;

    assign y0_2 = (x4_1 & x1_2) ^ (x4_2 & x1_1) ^ (x4_2 & x1_2) ^ x3_1 ^ (x2_1 & x1_1) ^ (x2_1 & x1_2) ^ (x2_2 & x1_1) ^ (x2_2 & x1_2) ^ (x1_1 & x0_1) ^ (x1_1 & x0_2) ^ (x1_2 & x0_1) ^ x1_2 ^ x0_2 ;
    assign y1_2 = x4_2 ^ (x3_0 & x2_2) ^ (x3_0 & x1_2) ^ (x3_2 & x2_0) ^ (x3_2 & x2_2) ^ (x3_2 & x1_0) ^ (x2_0 & x1_0) ^ (x2_0 & x1_2) ^ x2_0 ^ (x2_2 & x1_0) ^ x2_2 ^ x1_0 ^ x1_2 ;
    assign y2_2 = (x4_0 & x3_1) ^ (x4_1 & x3_0) ^ x2_0 ^ x1_1 ^ 1 ;
    assign y3_2 = (x4_0 & x0_2) ^ (x4_2 & x0_0) ^ (x4_2 & x0_2) ^ (x3_0 & x0_2) ^ (x3_2 & x0_0) ^ x3_2 ^ x2_2 ^ x1_0 ^ x0_0 ^ x0_2 ;
    assign y4_2 = (x4_0 & x1_0) ^ (x4_0 & x1_2) ^ (x4_2 & x1_0) ^ (x4_2 & x1_2) ^ x4_2 ^ x3_0 ^ x3_2 ^ (x1_0 & x0_2) ^ (x1_2 & x0_0) ^ (x1_2 & x0_2) ;    

endmodule
